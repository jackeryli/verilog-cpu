module mov (In1, In2);
input [31:0] In2;
output [31:0] In1;
assign In1 = In2;
endmodule