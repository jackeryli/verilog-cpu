module mov (In, Out);
input [31:0] In;
output [31:0] Out;
assign Out = In;
endmodule