module pc (count);
inout [7:0] count;
assign count = count+1;
endmodule
