module mov (In, Out);
input [31:0] In;
output wire [31:0] Out;
assign Out = In;
endmodule
